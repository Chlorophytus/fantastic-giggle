`timescale 1ns / 1ps
// Control Unit
module control
   (input wire logic aclk,
    input wire logic aresetn,

    // Enable this block
    input wire logic rx_enable);
endmodule: control
