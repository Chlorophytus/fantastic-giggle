../rtl_brancher/brancher.sv