`timescale 1ns / 1ps
module control_dut
   (input wire aclk,
    input wire aresetn,
    input wire rx_enable);

    control d(.*); 
endmodule
