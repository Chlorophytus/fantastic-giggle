../rtl_adder2/adder2.sv