../rtl_alu2/alu2.sv