../rtl_memory/memory.sv